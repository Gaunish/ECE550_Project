right_shift(input[31:0] operandA, 
			  input[4:0] shiftamt, 
			  output[31:0] result);
			  
endmodule